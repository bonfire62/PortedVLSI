`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    15:29:08 12/11/2017 
// Design Name: 
// Module Name:    Spiral_Rom 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Spiral_Rom(rom_row, col,  bit_out);
   input [6:0]rom_row;
   input [7:0]col;
   output bit_out;
   
   reg 	  [159:0]ROW;

   	always@(rom_row)
		case(rom_row)
			7'h0 : ROW = 120'b011111111111111110000000000000000000000000000011111111111111111111111111111111100000000000000000000000000000111111111111;
			7'h1 : ROW = 120'b111111111111100000000000000000000000011111111111111111111111111111111111111111111111111100000000000000000000000011111111;
			7'h2 : ROW = 120'b111111111100000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000011111;
			7'h3 : ROW = 120'b111111100000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000001;
			7'h4 : ROW = 120'b111000000000000000000111111111111111111111111111000000000000000000000000000001111111111111111111111111110000000000000000;
			7'h5 : ROW = 120'b100000000000000001111111111111111111111000000000000000000000000000000000000000000000001111111111111111111111000000000000;
			7'h6 : ROW = 120'b000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000001111111111111111111100000000;
			7'h7 : ROW = 120'b000000000011111111111111111000000000000000000000000000000000000000000000000000000000000000000000001111111111111111100000;
			7'h8 : ROW = 120'b000000011111111111111110000000000000000000000000000000001111111111111000000000000000000000000000000000111111111111111100;
			7'h9 : ROW = 120'b000011111111111111100000000000000000000000001111111111111111111111111111111111111000000000000000000000000011111111111111;
			7'hA : ROW = 120'b011111111111111100000000000000000000111111111111111111111111111111111111111111111111111110000000000000000000011111111111;
			7'hB : ROW = 120'b111111111111100000000000000000011111111111111111111111111111111111111111111111111111111111111100000000000000000001111111;
			7'hC : ROW = 120'b111111111100000000000000000111111111111111111111111111111111111111111111111111111111111111111111110000000000000000001111;
			7'hD : ROW = 120'b111111100000000000000001111111111111111111111100000000000000000000000000000000011111111111111111111111000000000000000011;
			7'hE : ROW = 120'b111100000000000000011111111111111111111000000000000000000000000000000000000000000000001111111111111111111100000000000000;
			7'hF : ROW = 120'b110000000000000011111111111111111000000000000000000000000000000000000000000000000000000000001111111111111111100000000000;
			7'h10 : ROW = 120'b000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000;
			7'h11 : ROW = 120'b000000000001111111111111100000000000000000000000000111111111111111111111110000000000000000000000000011111111111111100000;
			7'h12 : ROW = 120'b000000001111111111111100000000000000000000011111111111111111111111111111111111111100000000000000000000011111111111111000;
			7'h13 : ROW = 120'b000000111111111111100000000000000000011111111111111111111111111111111111111111111111111100000000000000000011111111111111;
			7'h14 : ROW = 120'b000011111111111100000000000000001111111111111111111111111111111111111111111111111111111111111000000000000000011111111111;
			7'h15 : ROW = 120'b001111111111100000000000000001111111111111111111111111000000000000000011111111111111111111111111000000000000000011111111;
			7'h16 : ROW = 120'b111111111110000000000000011111111111111111111000000000000000000000000000000000001111111111111111111100000000000000111111;
			7'h17 : ROW = 120'b111111111000000000000011111111111111111000000000000000000000000000000000000000000000001111111111111111100000000000000111;
			7'h18 : ROW = 120'b111111100000000000001111111111111110000000000000000000000000000000000000000000000000000000111111111111111100000000000001;
			7'h19 : ROW = 120'b111110000000000001111111111111100000000000000000000000000000000000000000000000000000000000000011111111111111000000000000;
			7'h1A : ROW = 120'b111000000000000111111111111100000000000000000000011111111111111111111111111100000000000000000000011111111111111000000000;
			7'h1B : ROW = 120'b100000000000011111111111100000000000000000011111111111111111111111111111111111111100000000000000000011111111111110000000;
			7'h1C : ROW = 120'b000000000001111111111100000000000000001111111111111111111111111111111111111111111111111000000000000000011111111111100000;
			7'h1D : ROW = 120'b000000000111111111110000000000000011111111111111111111111111111111111111111111111111111111100000000000000111111111111000;
			7'h1E : ROW = 120'b000000011111111111000000000000011111111111111111111100000000000000000000011111111111111111111100000000000001111111111100;
			7'h1F : ROW = 120'b000000111111111100000000000011111111111111111000000000000000000000000000000000001111111111111111100000000000001111111111;
			7'h20 : ROW = 120'b000011111111110000000000001111111111111100000000000000000000000000000000000000000000011111111111111000000000000111111111;
			7'h21 : ROW = 120'b000111111111000000000000111111111111100000000000000000000000000000000000000000000000000011111111111110000000000001111111;
			7'h22 : ROW = 120'b011111111110000000000011111111111100000000000000000000001111111111111000000000000000000000011111111111110000000000011111;
			7'h23 : ROW = 120'b111111111000000000001111111111100000000000000000011111111111111111111111111100000000000000000011111111111000000000001111;
			7'h24 : ROW = 120'b111111110000000000111111111110000000000000001111111111111111111111111111111111111000000000000000111111111110000000000011;
			7'h25 : ROW = 120'b111111100000000001111111111000000000000011111111111111111111111111111111111111111111100000000000001111111111100000000001;
			7'h26 : ROW = 120'b111110000000000111111111100000000000001111111111111111111111000001111111111111111111111100000000000011111111110000000000;
			7'h27 : ROW = 120'b111100000000001111111110000000000001111111111111111000000000000000000000001111111111111111000000000000111111111100000000;
			7'h28 : ROW = 120'b111000000000011111111100000000000111111111111100000000000000000000000000000000011111111111110000000000001111111110000000;
			7'h29 : ROW = 120'b110000000001111111110000000000011111111111100000000000000000000000000000000000000011111111111100000000000111111111000000;
			7'h2A : ROW = 120'b100000000011111111100000000001111111111100000000000000000000000000000000000000000000011111111111000000000001111111110000;
			7'h2B : ROW = 120'b100000000111111111000000000011111111110000000000000000111111111111111110000000000000000111111111110000000000111111111000;
			7'h2C : ROW = 120'b000000001111111110000000001111111111000000000000001111111111111111111111111000000000000001111111111000000000011111111100;
			7'h2D : ROW = 120'b000000001111111100000000011111111100000000000001111111111111111111111111111111100000000000011111111110000000001111111100;
			7'h2E : ROW = 120'b000000011111111000000000111111111000000000001111111111111111111111111111111111111000000000000111111111000000000111111110;
			7'h2F : ROW = 120'b000000111111110000000001111111110000000000111111111111111000000000001111111111111110000000000011111111100000000011111111;
			7'h30 : ROW = 120'b000000111111100000000011111111100000000011111111111100000000000000000000011111111111100000000001111111110000000001111111;
			7'h31 : ROW = 120'b000001111111100000000111111111000000000111111111100000000000000000000000000011111111111000000000111111111000000001111111;
			7'h32 : ROW = 120'b000001111111000000000111111110000000001111111110000000000000000000000000000000111111111100000000011111111100000000111111;
			7'h33 : ROW = 120'b000011111111000000001111111100000000011111111000000000000000000000000000000000001111111110000000001111111100000000011111;
			7'h34 : ROW = 120'b000011111110000000011111111000000000111111110000000000011111111111111100000000000011111111000000000111111110000000011111;
			7'h35 : ROW = 120'b000111111110000000011111111000000001111111100000000001111111111111111111000000000001111111100000000011111111000000001111;
			7'h36 : ROW = 120'b000111111110000000011111110000000011111111000000000111111111111111111111110000000000111111110000000011111111000000001111;
			7'h37 : ROW = 120'b000111111100000000111111110000000011111111000000001111111111111111111111111100000000011111111000000001111111100000000111;
			7'h38 : ROW = 120'b000111111100000000111111110000000011111110000000011111111100000000011111111110000000011111111000000001111111100000000111;
			7'h39 : ROW = 120'b000111111100000000111111100000000111111110000000011111110000000000000111111111000000001111111100000000111111100000000111;
			7'h3A : ROW = 120'b000111111100000000111111100000000111111110000000011111110000000000000011111111000000001111111100000000111111100000000111;
			7'h3B : ROW = 120'b000111111100000000111111100000000111111110000000011111110000010000000001111111100000000111111100000000111111110000000111;
			7'h3C : ROW = 120'b000111111100000000111111110000000111111110000000011111111000111100000000111111100000000111111100000000111111110000000011;
			7'h3D : ROW = 120'b000111111100000000111111110000000011111110000000001111111111111100000000111111100000000111111100000000111111110000000011;
			7'h3E : ROW = 120'b000111111110000000011111110000000011111111000000000111111111111100000000111111100000000111111100000000111111110000000011;
			7'h3F : ROW = 120'b000111111110000000011111111000000001111111100000000001111111110000000001111111100000000111111100000000111111110000000111;
			7'h40 : ROW = 120'b000011111110000000011111111000000001111111110000000000000000000000000011111111000000001111111100000000111111100000000111;
			7'h41 : ROW = 120'b000011111111000000001111111100000000111111111000000000000000000000000111111111000000001111111100000000111111100000000111;
			7'h42 : ROW = 120'b000011111111000000001111111100000000011111111110000000000000000000001111111110000000011111111000000001111111100000000111;
			7'h43 : ROW = 120'b000001111111100000000111111110000000000111111111100000000000000001111111111100000000011111111000000001111111000000000111;
			7'h44 : ROW = 120'b000001111111100000000011111111000000000011111111111111000000011111111111110000000000111111110000000011111111000000001111;
			7'h45 : ROW = 120'b000000111111110000000001111111100000000000111111111111111111111111111111100000000001111111100000000011111111000000001111;
			7'h46 : ROW = 120'b000000011111111000000000111111111000000000001111111111111111111111111110000000000011111111000000000111111110000000011111;
			7'h47 : ROW = 120'b000000011111111100000000011111111100000000000001111111111111111111110000000000001111111110000000001111111100000000011111;
			7'h48 : ROW = 120'b000000001111111110000000001111111111000000000000000111111111111100000000000000011111111100000000011111111100000000111111;
			7'h49 : ROW = 120'b000000000111111111000000000111111111110000000000000000000000000000000000000001111111111000000000111111111000000001111111;
			7'h4A : ROW = 120'b100000000011111111100000000001111111111110000000000000000000000000000000001111111111100000000001111111110000000001111111;
			7'h4B : ROW = 120'b110000000001111111110000000000011111111111110000000000000000000000000001111111111111000000000011111111100000000011111111;
			7'h4C : ROW = 120'b111000000000111111111100000000000111111111111111000000000000000000011111111111111100000000000111111111000000000111111110;
			7'h4D : ROW = 120'b111100000000001111111110000000000001111111111111111111111111111111111111111111110000000000011111111110000000001111111100;
			7'h4E : ROW = 120'b111110000000000111111111100000000000001111111111111111111111111111111111111110000000000000111111111000000000011111111100;
			7'h4F : ROW = 120'b111111000000000011111111111000000000000001111111111111111111111111111111110000000000000011111111110000000000111111111000;
			7'h50 : ROW = 120'b111111110000000000111111111110000000000000000011111111111111111111111000000000000000001111111111100000000001111111110000;
			7'h51 : ROW = 120'b111111111000000000001111111111110000000000000000000000011111100000000000000000000001111111111110000000000111111111000000;
			7'h52 : ROW = 120'b011111111110000000000011111111111100000000000000000000000000000000000000000000001111111111111000000000001111111110000000;
			7'h53 : ROW = 120'b001111111111000000000000111111111111110000000000000000000000000000000000000001111111111111100000000000111111111100000000;
			7'h54 : ROW = 120'b000011111111110000000000001111111111111111000000000000000000000000000000011111111111111110000000000001111111111000000000;
			7'h55 : ROW = 120'b000001111111111100000000000001111111111111111111100000000000000000111111111111111111110000000000000111111111100000000001;
			7'h56 : ROW = 120'b000000011111111111000000000000001111111111111111111111111111111111111111111111111110000000000000011111111111000000000011;
			7'h57 : ROW = 120'b000000000111111111110000000000000001111111111111111111111111111111111111111111110000000000000001111111111100000000001111;
			7'h58 : ROW = 120'b000000000001111111111110000000000000000011111111111111111111111111111111111000000000000000001111111111110000000000011111;
			7'h59 : ROW = 120'b100000000000011111111111100000000000000000000011111111111111111111111000000000000000000000111111111111000000000001111111;
			7'h5A : ROW = 120'b111000000000000111111111111100000000000000000000000000000000000000000000000000000000000111111111111100000000000011111111;
			7'h5B : ROW = 120'b111110000000000001111111111111110000000000000000000000000000000000000000000000000001111111111111110000000000001111111111;
			7'h5C : ROW = 120'b111111100000000000001111111111111111000000000000000000000000000000000000000000011111111111111110000000000000111111111110;
			7'h5D : ROW = 120'b111111111000000000000001111111111111111111000000000000000000000000000000011111111111111111110000000000000011111111111000;
			7'h5E : ROW = 120'b111111111110000000000000001111111111111111111111111111000000011111111111111111111111111110000000000000001111111111100000;
			7'h5F : ROW = 120'b011111111111110000000000000000111111111111111111111111111111111111111111111111111111100000000000000001111111111110000000;
			7'h60 : ROW = 120'b000011111111111100000000000000000011111111111111111111111111111111111111111111111000000000000000000111111111111000000000;
			7'h61 : ROW = 120'b000000111111111111100000000000000000000011111111111111111111111111111111111000000000000000000000111111111111100000000000;
			7'h62 : ROW = 120'b000000001111111111111110000000000000000000000000011111111111111111000000000000000000000000001111111111111110000000000001;
			7'h63 : ROW = 120'b000000000001111111111111110000000000000000000000000000000000000000000000000000000000000001111111111111110000000000000111;
			7'h64 : ROW = 120'b000000000000001111111111111111100000000000000000000000000000000000000000000000000000111111111111111110000000000000011111;
			7'h65 : ROW = 120'b110000000000000001111111111111111111000000000000000000000000000000000000000000011111111111111111110000000000000001111111;
			7'h66 : ROW = 120'b111110000000000000001111111111111111111111100000000000000000000000000000111111111111111111111110000000000000001111111111;
			7'h67 : ROW = 120'b111111100000000000000000111111111111111111111111111111111111111111111111111111111111111111100000000000000000111111111111;
			7'h68 : ROW = 120'b111111111100000000000000000011111111111111111111111111111111111111111111111111111111111000000000000000000111111111111100;
			7'h69 : ROW = 120'b111111111111100000000000000000000011111111111111111111111111111111111111111111111000000000000000000000111111111111110000;
			7'h6A : ROW = 120'b001111111111111110000000000000000000000001111111111111111111111111111111110000000000000000000000001111111111111110000000;
			7'h6B : ROW = 120'b000001111111111111110000000000000000000000000000000000000000000000000000000000000000000000000001111111111111110000000000;
			7'h6C : ROW = 120'b000000011111111111111111100000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000;
			7'h6D : ROW = 120'b000000000001111111111111111111000000000000000000000000000000000000000000000000000000011111111111111111110000000000000001;
			7'h6E : ROW = 120'b000000000000001111111111111111111111000000000000000000000000000000000000000000011111111111111111111110000000000000000111;
			7'h6F : ROW = 120'b100000000000000000111111111111111111111111111100000000000000000000000111111111111111111111111111100000000000000000111111;
			7'h70 : ROW = 120'b111100000000000000000001111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111111111;
			7'h71 : ROW = 120'b111111100000000000000000000011111111111111111111111111111111111111111111111111111111111000000000000000000000111111111111;
			7'h72 : ROW = 120'b111111111110000000000000000000000011111111111111111111111111111111111111111111111000000000000000000000001111111111111110;
			7'h73 : ROW = 120'b111111111111111000000000000000000000000000001111111111111111111111111110000000000000000000000000000011111111111111110000;
			7'h74 : ROW = 120'b011111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000;
			7'h75 : ROW = 120'b000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000;
			7'h76 : ROW = 120'b000000000111111111111111111111000000000000000000000000000000000000000000000000000000011111111111111111111100000000000000;
			7'h77 : ROW = 120'b000000000000111111111111111111111111110000000000000000000000000000000000000001111111111111111111111111100000000000000000;
			default: ROW = 120'b000000000000111111111111111111111111110000000000000000000000000000000000000001111111111111111111111111100000000000000000;

		endcase
		
		assign bit_out = ROW[col];

endmodule
